module MTran_Lab1_Verilog_AndGate(a,b,y);

input a,b;
output y;
and (y,a,b);

endmodule